module lab1part1 ();

// Check to see if other modules work --> DFF, MUX, and counter

endmodule
